`include "lift_controller.sv"
`include "lift_trans.sv"
`include "lift_gen.sv"
`include "lift_intf.sv"
`include "lift_bfm.sv"
`include "lift_env.sv"
`include "lift_test.sv"
`include "lift_controller_tb.sv"





